VCF

Vin 1 0 AC 50m

Xstage1 1 2 3 0 stage
Xstage2 2 3 4 0 stage
Xstage3 3 4 5 0 stage
Xstage4 4 5 0 0 stage

.subckt stage 3 8 12 0
VDD 1 0 DC 2.5
VSS 2 0 DC -2.5

Vabc 4 0 DC 2.5

R1 3 6 100K
R2 6 0 220

C1 7 12 100pico

R3 8 9 100K
R4 9 0 200

R5 8 2 10K

Rabc 4 10 20K

*        Amplifier Bias Input
*        |  Diode Bias
*        |  | Positive Input
*        |  | | Negative Input
*        |  | | | Output
*        |  | | | | Negative power supply
*        |  | | | | | Buffer Input
*        |  | | | | | | Buffer Output
*        |  | | | | | | | Positive power supply
*        |  | | | | | | | |
Xopamp1 10 11 6 9 7 2 7 8 1 LM13700/NS
.ends
*.ac dec 10000 1Hz 50kHz
*.tran 1u 10m
*.plot V(3) V(5) V(8)
*.op

* \\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\            
* LM13700 Dual Operational Transconductance Amplifier                 
* \\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\                 
*
*                  Amplifier Bias Input
*                  | Diode Bias
*                  | | Positive Input
*                  | | | Negative Input
*                  | | | | Output
*                  | | | | | Negative power supply
*                  | | | | | | Buffer Input
*                  | | | | | | | Buffer Output
*                  | | | | | | | | Positive power supply
*                  | | | | | | | | |
.subckt LM13700/NS 1 2 3 4 5 6 7 8 11
	*
	* Features:
	* gm adjustable over 6 decades.
	* Excellent gm linearity.
	* Linearizing diodes.
	* Wide supply range of +/-2V to +/-22V.
	*
	* Note:  This model is single-pole in nature and over-estimates
	*       AC bandwidth and phase margin (stability) by over 2X.   
	*       Although refinement may be possible in the future, please
	*       use benchtesting to finalize AC circuit design.
	* 
	* Note: Model is for single device only and simulated
	*       supply current is 1/2 of total device current.
	*
	******************************************************
	* 
	C1  6  4  4.8P
	C2  3  6  4.8P
	* Output capacitor  
	C3  5  6  6.26P                                       
	D1  2  4  DX
	D2  2  3  DX
	D3  11 21 DX
	D4  21 22 DX
	D5  1  26 DX
	D6  26 27 DX
	D7  5  29 DX
	D8  28 5  DX
	D10 31 25 DX
	* Clamp for -CMR  
	D11 28 25 DX                                        
	* Ios source 
	F1  4  3  POLY(1)   V6 1E-10 5.129E-2 -1.189E4 1.123E9 
	F2  11 5  V2        1.022
	F3  25 6  V3        1.0
	F4  5  6  V1        1.022
	* Output impedance 
	F5  5  0  POLY(2)   V3 V7 0 0 0 0 1                  
	G1  0  33 5         0 .55E-3
	I1  11 6  300U
	Q1  24 32 31        QX1
	Q2  23 3  31        QX2
	Q3  11 7  30        QZ
	Q4  11 30 8         QY
	V1  22 24 0V
	V2  22 23 0V
	V3  27 6  0V
	V4  11 29 1.4
	V5  28 6  1.2
	V6  4  32 0V
	V7  33 0  0V
	.model QX1 NPN (IS=5E-16     BF=200 NE=1.15 ISE=.63E-16 IKF=1E-2)
	.model QX2 NPN (IS=5.125E-16 BF=200 NE=1.15 ISE=.63E-16 IKF=1E-2)
	.model QY  NPN (IS=6E-15     BF=50)
	.model QZ  NPN (IS=5E-16     BF=266)  
	.model DX  D   (IS=5E-16)
.ends

.end
